module lorentz();

reg [63:0] a,b,c;


initial
begin
	a = 64'h4024000000000000; //a = 10
	b = 64'h403C000000000000' //b = 28
	c = 64'h4005555555555555; // c = 8/3
end